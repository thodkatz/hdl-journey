module main;
  initial
    begin
      $display("Hello Verilog");
      $finish;
    end
endmodule
